interface spi_if #(parameter CLK_DIV = 4)(
     input logic clk, 
     input logic rst_n
);

    // DUT interface signals
    logic        start;
    logic [7:0]  tx_data;
    logic [7:0]  rx_data;
    logic        busy;
    logic        done;

    // SPI physical interface
    logic        sclk;
    logic        mosi;
    logic        miso;
    logic        cs_n;

    // Clocking block for driver
    clocking drv_cb @(posedge clk);
        default input #1ns output #1ns;
        output start, tx_data;
        input  busy, done, rx_data;
        output mosi, cs_n, sclk;
        input  miso;
    endclocking

    // Clocking block for monitor
    clocking mon_cb @(posedge clk);
        default input #1ns output #1ns;
        input start, tx_data, busy, done, rx_data;
        input mosi, cs_n, sclk, miso;
    endclocking

    // Modports for separation of roles
    modport drv_mp  (clocking drv_cb);
    modport mon_mp (clocking mon_cb);

endinterface
