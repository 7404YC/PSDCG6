// T013: Ensure MOSI only changes on rising sclk edges
property T013;
	@(posedge clk)
	disable iff (!rst_n)
		(
			// When there is no rising sclk events, but detect mosi changes, this will flag error
			!($rose(sclk)) |-> (mosi === $past(mosi))
		);
endproperty
ASSERT_T013: assert property (T013)
	else $error("ASSERT ", $sformatf("Error T013"));

// T018: When the SPI is idle, ensure no sclk events and cs_n is pulled high.
property T018;
	@(posedge clk)
	disable iff (!rst_n)
		(
			(state == 0 && start == 0) |->
			(
				sclk == 0 &&
				cs_n == 1
			)
		);
endproperty
ASSERT_T018: assert property (T018)
	else $error("ASSERT ", $sformatf("Error T018"));

// T020: All outputs are set to default/reset values when rst_n = 0, except mosi
// Reason to use always_comb is because the reset is asynchronous to the clock, so we cannot use property which is sensitive to the clock
always_comb begin
	if (rst_n == 1'b0) begin
	ASSERT_T020:
		assert final (
					(busy == 1'b0) &&
					(done == 1'b0) &&
					(rx_data == 8'b0) &&
					(sclk == 1'b0) &&
					(cs_n == 1'b1)
				)
		else $error("ASSERT ", $sformatf("Error T020"));
	end
end

// T025: Ensure no glitch on sclk rising edge
property T025;
	@(posedge clk)
	disable iff (!rst_n || !busy)
	$rose(sclk) |-> ##1 (sclk == 1) ##(CLK_DIV/2-1) $fell(sclk);
endproperty
ASSERT_T025:
	assert property (T025)
	else $error ("ASSERT ", $sformatf("Error T025"));

// T026: Ensure no glitch on sclk falling edge
property T026;
	@(posedge clk)
	disable iff (!rst_n || !busy)
	$fell(sclk) |-> ##1 (sclk == 0) ##(CLK_DIV/2-1) $rose(sclk);
endproperty
ASESRT_T026:
	assert property (T026)
	else $error ("ASSERT ", $sformatf("Error T026"));


